// ATS Library 
// Library contains 
// - Processor Defines 
// 
//==============================================================

// RISCV Processor Defines 
`define RV_IMEM_WIDTH 32
`define RV_IMEM_DEPTH 256
`define RV_DMEM_WIDTH 32
`define RV_DMEM_DEPTH 256       // 256
`define RV_RF_WIDTH 32          // Register File Wdith
`define RV_RF_DEPTH 32          // Register File Depth

